package apb_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "apb_packet.sv"
`include "apb_monitor.sv"
`include "apb_sequencer.sv"
`include "apb_seq.sv"
`include "apb_master_driver.sv"
`include "apb_slave_driver.sv"
`include "apb_agent.sv"


endpackage: apb_pkg
